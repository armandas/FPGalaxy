library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity explosion_rom is
    port(
        addr: in std_logic_vector(9 downto 0);
        data: out std_logic_vector(2 downto 0)
    );
end explosion_rom;

architecture content of explosion_rom is
    type rgb_array is array(0 to 31) of std_logic_vector(2 downto 0);
    type rom_type is array(0 to 31) of rgb_array;

    signal rgb_row: rgb_array;

    constant EXPLOSION: rom_type :=
    (
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "111", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "110", "111", "110", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "111", "111", "000", "000", "100", "000", "000", "000", "100", "000", "111", "110", "110", "110", "000", "000", "100", "100", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "111", "110", "110", "110", "111", "000", "000", "100", "000", "110", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "111", "110", "110", "110", "110", "111", "100", "100", "111", "111", "110", "100", "110", "111", "111", "000", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "100", "000", "111", "110", "110", "100", "110", "110", "110", "110", "110", "110", "100", "110", "110", "111", "111", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "111", "110", "100", "100", "100", "110", "100", "100", "100", "100", "100", "100", "110", "110", "110", "110", "110", "110", "110", "111", "111", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "100", "000", "111", "111", "110", "100", "100", "110", "110", "000", "110", "100", "110", "100", "100", "100", "100", "110", "110", "111", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "110", "000", "100", "100", "110", "000", "000", "000", "000", "100", "100", "110", "110", "111", "111", "110", "110", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "100", "000", "111", "111", "000", "110", "110", "000", "100", "100", "100", "100", "100", "000", "000", "110", "111", "111", "000", "000", "000", "100", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "111", "111", "111", "111", "110", "110", "110", "100", "000", "110", "110", "100", "000", "100", "100", "100", "000", "000", "000", "000", "100", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "111", "111", "110", "110", "110", "100", "000", "100", "110", "100", "100", "000", "110", "110", "110", "100", "110", "100", "111", "111", "111", "111", "111", "111", "111", "000", "000", "000"),
        ("000", "000", "000", "111", "111", "110", "110", "100", "100", "000", "110", "110", "100", "100", "100", "110", "100", "100", "110", "000", "110", "110", "100", "110", "110", "110", "100", "110", "111", "000", "000", "000"),
        ("000", "000", "000", "000", "111", "111", "111", "110", "110", "000", "100", "100", "100", "100", "110", "110", "000", "100", "100", "100", "100", "100", "100", "100", "100", "100", "100", "110", "111", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "100", "111", "111", "111", "110", "110", "110", "100", "000", "000", "100", "100", "000", "110", "100", "110", "110", "000", "110", "110", "100", "100", "110", "111", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "100", "000", "111", "111", "110", "110", "100", "110", "110", "100", "100", "110", "100", "000", "111", "111", "111", "111", "110", "110", "110", "111", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "110", "100", "000", "000", "111", "110", "000", "100", "110", "110", "000", "110", "110", "100", "100", "110", "111", "111", "111", "111", "111", "111", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "111", "110", "110", "100", "000", "110", "100", "100", "100", "110", "110", "100", "110", "110", "111", "111", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "110", "000", "000", "111", "110", "100", "100", "110", "110", "100", "100", "110", "100", "000", "100", "100", "000", "110", "111", "111", "100", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "111", "110", "100", "100", "110", "000", "000", "110", "110", "110", "110", "000", "000", "100", "100", "100", "110", "100", "111", "110", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "100", "000", "111", "000", "000", "110", "000", "100", "100", "100", "100", "100", "100", "111", "110", "000", "110", "110", "100", "110", "111", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "100", "111", "111", "110", "100", "100", "100", "100", "100", "000", "110", "100", "100", "111", "111", "111", "111", "110", "110", "100", "111", "111", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "111", "110", "100", "100", "110", "110", "110", "100", "100", "110", "100", "110", "111", "000", "000", "000", "111", "111", "111", "110", "111", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "110", "100", "111", "110", "100", "110", "000", "100", "100", "100", "110", "110", "110", "100", "111", "000", "110", "000", "100", "000", "000", "111", "111", "111", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "111", "110", "100", "110", "110", "110", "110", "100", "000", "100", "100", "000", "111", "100", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "100", "000", "000", "111", "111", "111", "111", "111", "111", "111", "111", "110", "100", "100", "110", "111", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "111", "111", "111", "100", "000", "000", "000", "000", "111", "111", "110", "110", "110", "111", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "110", "000", "100", "000", "000", "111", "111", "111", "111", "111", "000", "100", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000"),
        ("000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000", "000")
    );
begin
    rgb_row <= EXPLOSION(conv_integer(addr(9 downto 5)));
    data <= rgb_row(conv_integer(addr(4 downto 0)));
end content;
